module core_top(
    input wire clk,
    input wire reset
);

// To Implement

endmodule
